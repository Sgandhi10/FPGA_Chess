module DD2_Final_PRJ ();
	
endmodule